/*
 * ame_ver_mem.sv
 *
 *  Created on: 2022-07-16 22:07
 *      Author: Jack Chen <redchenjs@live.com>
 */

`timescale 1 ns / 1 ps

module ame_ver_mem(
    input logic clk_i,
    input logic rst_n_i,

    output logic ame_run,
    output logic ame_done,
    output logic ame_error
);

endmodule
